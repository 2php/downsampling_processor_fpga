module test1mem ()

endmodule