
module unnamed (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
